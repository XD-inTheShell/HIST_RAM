module SRAM_SC_s10_user_rst_clkgate_2 (
		output wire  ninit_done  // ninit_done.ninit_done
	);
endmodule

