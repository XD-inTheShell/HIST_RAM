module SRAM_SC_iopll_0 (
		input  wire  rst,      //   reset.reset
		input  wire  refclk,   //  refclk.clk
		output wire  locked,   //  locked.export
		output wire  outclk_0  // outclk0.clk
	);
endmodule

