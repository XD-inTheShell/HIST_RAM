module SRAM_SC_clock_bridge_0 (
		input  wire  in_clk,  //  in_clk.clk
		output wire  out_clk  // out_clk.clk
	);
endmodule

