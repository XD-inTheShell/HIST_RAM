module SRAM_SC_reset_in (
		input  wire  in_reset,  //  in_reset.reset
		output wire  out_reset  // out_reset.reset
	);
endmodule

